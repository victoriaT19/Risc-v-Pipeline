`timescale 1ns / 1ps

module Controller (
    //Input
    input logic [6:0] Opcode,
    //7-bit opcode field from the instruction

    //Outputs
    output logic ALUSrc,
    //0: The second ALU operand comes from the second register file output (Read data 2); 
    //1: The second ALU operand is the sign-extended, lower 16 bits of the instruction.
    output logic MemtoReg,
    //0: The value fed to the register Write data input comes from the ALU.
    //1: The value fed to the register Write data input comes from the data memory.
    output logic RegWrite, //The register on the Write register input is written with the value on the Write data input 
    output logic MemRead,  //Data memory contents designated by the address input are put on the Read data output
    output logic MemWrite, //Data memory contents designated by the address input are replaced by the value on the Write data input.
    output logic [1:0] ALUOp,  //00: LW/SW; 01:Branch; 10: Rtype; 11: JAL
    output logic Branch,  //0: branch is not taken; 1: branch is taken
    output logic JalrSel, // flag para Jalr
    output logic Halt,
    output logic RWSel
);

  logic [6:0] R_TYPE, I_TYPE, LW, SW, BR, JAL, JALR, HALT; //adicionado as instruc�es do tipo I, JAL e JALR e pseudo-instru��o HALT

  assign R_TYPE = 7'b0110011;  //add, sub, and, xor, or, slt
  assign I_TYPE = 7'b0010011; //addi, slti, slli, srli, srai
  assign LW = 7'b0000011;  //lw, lb, lh, lbu
  assign SW = 7'b0100011;  //sw, sb, sh
  assign BR = 7'b1100011;  //beq, bne, blt, bge
  assign JAL = 7'b1101111; //adicionado o opcode da instruc�o jal
  assign JALR = 7'b1100111; //adicionado o opcode da instruc�o jalr
  assign HALT = 7'b1111111; /*-> opcode inventado*/

  assign ALUSrc = (Opcode == LW || Opcode == SW || Opcode == I_TYPE || Opcode == JALR); //adicionado as instruc�es do tipo I e JALR
  assign MemtoReg = (Opcode == LW);
  assign RegWrite = (Opcode == R_TYPE || Opcode == LW || Opcode == I_TYPE || Opcode == JAL || Opcode == JALR); //adicionado as instruc�es do tipo I, JAL e JALR
  assign MemRead = (Opcode == LW);
  assign MemWrite = (Opcode == SW);
  assign ALUOp[0] = (Opcode == BR || Opcode == JAL);
  assign ALUOp[1] = (Opcode == R_TYPE || Opcode == I_TYPE || Opcode == JAL); 
  assign Branch = (Opcode == BR || Opcode == JAL);
  assign JalrSel = (Opcode == JALR); 
  assign Halt = (Opcode == HALT);
  assign RWSel = (Opcode == JAL || Opcode == JALR);
  
endmodule